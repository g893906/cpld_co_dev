/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ*********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   led������ʵ��
**********************************************************************/

module led1(led);
	output[7:0] led;
	  assign led=8'b00000000; //����ȫ��8��led
	//  assign led=8'b01010101;//�Զ��led����
                          //ʹ��������ֵ���assignʵ��
endmodule


