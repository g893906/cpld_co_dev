/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   ���뿪����������LED
********************************************************************/


module ckey_led(ckey,led);
  input  [4:1] ckey;                   // ckey[1]  ~ ckey[4]
  output [4:1] led;                    // led[1] ~ led[4]
   

// ��������led[1]����led[8]���ң���1����0��
// ��������ckey��Ϊ0���ر�Ϊ1
assign led = ckey;

endmodule