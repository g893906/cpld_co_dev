/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   led����˸ʵ��
********************************************************************/




module led_twinkle(led,clk);// ģ�������˿ڲ���
	output [8:1] led;
	input clk;
	reg[8:1] led;// ����˿ڶ���Ϊ�Ĵ�����
	reg[24:0] counter;  // �м����counter����Ϊ�Ĵ�����
	
	always@(posedge clk)//��ʱ�Ӹ�������
		begin // ˳����䣬��endֹ
			counter<=counter+1;  //<=�� =����
		    //if(counter==25'b1011111010111100001000000) //�б�counter�е���ֵΪ25000000ʱ
		    if(counter==25'd25000000)
			
				begin	
					led<=~led;// led[1]-led[8]��תһ��
			 		counter<=0;//���¼���
				end   
		end
endmodule
	