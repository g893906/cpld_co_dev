/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   ��ȡ�����ź�ʵ��
********************************************************************/


module key_led(key,led);//
input[6:1]key;
output[6:1]led;
reg[6:1]led_r;
reg[6:1]buffer;
assign led=led_r;

always@(key)
begin
	buffer=key;
	case(buffer)
		6'b111110:led_r=6'b111110;//������µ���key1,��ô����LED1
		6'b111101:led_r=6'b111100;//������µ���key2,��ô����LED1-LED2
		6'b111011:led_r=6'b111000;//key3
		6'b110111:led_r=6'b110000;//key4
	   6'b101111:led_r=6'b100000;//key5
	   6'b011111:led_r=6'b000000;//key6
	    
		default:led_r=6'b111111;
	endcase
end
endmodule